
  `timescale 1ns/1ps
//==============================================================================
//
//
//
//
//
//
//
//
//==============================================================================

  module Test_Top (
  
    input    wire    sys_clk ,
    input    wire    sys_rst ,
    output   wire    data_o  
  
  );
//----------------------------

   assign data_o = 1'b0 ;


  endmodule
